-- This Source Code Form is subject to the terms of the Mozilla Public
-- License, v. 2.0. If a copy of the MPL was not distributed with this file,
-- You can obtain one at http://mozilla.org/MPL/2.0/.
--
-- Copyright (c) 2014-2026, Lars Asplund lars.anders.asplund@gmail.com

context com_context is
  library vunit_lib;

  use vunit_lib.codec_2008p_pkg.all;
  use vunit_lib.codec_builder_2008p_pkg.all;
  use vunit_lib.codec_builder_pkg.all;
  use vunit_lib.codec_pkg.all;
  use vunit_lib.com_common_pkg.all;
  use vunit_lib.com_debug_codec_builder_pkg.all;
  use vunit_lib.com_deprecated_pkg.all;
  use vunit_lib.com_pkg.all;
  use vunit_lib.com_string_pkg.all;
  use vunit_lib.com_types_pkg.all;
end context;
