library ieee;
use ieee.std_logic_1164.all;

architecture arch of buffer1 is

begin
    Q <= D;
end architecture;
