-- This Source Code Form is subject to the terms of the Mozilla Public
-- License, v. 2.0. If a copy of the MPL was not distributed with this file,
-- You can obtain one at http://mozilla.org/MPL/2.0/.
--
-- Copyright (c) 2014-2022, Lars Asplund lars.anders.asplund@gmail.com

context data_types_context is
  library vunit_lib;
  use vunit_lib.types_pkg.all;
  use vunit_lib.integer_vector_ptr_pkg.all;
  use vunit_lib.integer_vector_ptr_pool_pkg.all;
  use vunit_lib.integer_array_pkg.all;
  use vunit_lib.queue_pkg.all;
  use vunit_lib.queue_pool_pkg.all;
  use vunit_lib.string_ptr_pkg.all;
  use vunit_lib.string_ptr_pool_pkg.all;
  use vunit_lib.byte_vector_ptr_pkg.all;
  use vunit_lib.dict_pkg.all;
end context;
