-- This Source Code Form is subject to the terms of the Mozilla Public
-- License, v. 2.0. If a copy of the MPL was not distributed with this file,
-- You can obtain one at http://mozilla.org/MPL/2.0/.
--
-- Copyright (c) 2015-2016, Lars Asplund lars.anders.asplund@gmail.com

use std.env.stop;

package body vunit_stop_pkg is
  procedure vunit_stop(status : integer) is
  begin
    stop(status);
  end procedure;
end package body;
