// This Source Code Form is subject to the terms of the Mozilla Public
// License, v. 2.0. If a copy of the MPL was not distributed with this file,
// You can obtain one at http://mozilla.org/MPL/2.0/.
//
// Copyright (c) 2014-2015, Lars Asplund lars.anders.asplund@gmail.com

module simple();
   always begin
      #1;
      $display("hello");
      #1;
   end
endmodule
