-- This Source Code Form is subject to the terms of the Mozilla Public
-- License, v. 2.0. If a copy of the MPL was not distributed with this file,
-- You can obtain one at http://mozilla.org/MPL/2.0/.
--
-- Copyright (c) 2015, Lars Asplund lars.anders.asplund@gmail.com

package body vunit_stop_pkg is
  procedure vunit_stop(status : integer) is
  begin
    std.env.stop(status);
  end procedure;
end package body;
