library ieee;
use ieee.std_logic_1164.all;

entity buffer1 is
  port (
    D : in std_logic;
    Q : out std_logic
  );
end entity;
